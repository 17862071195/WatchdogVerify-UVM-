class c_4_3;
    rand integer delay; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq_lib/watchdog_resen_virtual_sequence.sv:21)
    {
       (delay inside {[5:3]});
    }
endclass

program p_4_3;
    c_4_3 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zzzzx0zxz1z0zz11xx01x1z110000zzzxzxzxxxxxxxxxxxzxzzxzzxxxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
