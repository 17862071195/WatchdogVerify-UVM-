class c_41_3;
    rand integer delay; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq_lib/watchdog_resen_virtual_sequence.sv:21)
    {
       (delay inside {[5:3]});
    }
endclass

program p_41_3;
    c_41_3 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x10z0z00z10z001zxx01x100zxxzz0zzzzzzxxzxzzzzxxxzxxxzzzzxzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
