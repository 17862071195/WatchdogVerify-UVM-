class c_46_3;
    rand integer delay; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq_lib/watchdog_resen_virtual_sequence.sv:21)
    {
       (delay inside {[5:3]});
    }
endclass

program p_46_3;
    c_46_3 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx000z01x0xz1z0zx0x1zxz01100zx0zzzzzxzxxxzzzxxzzxzzzxzzxzzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
