`ifndef WATCHDOG_TESTS_SVH
`define WATCHDOG_TESTS_SVH

	`include "watchdog_base_test.sv"
	`include "watchdog_integration_test.sv"
	`include "watchdog_regacc_test.sv"
	`include "watchdog_apbacc_test.sv"

	`include "watchdog_countdown_test.sv"
	`include "watchdog_reload_test.sv"
	`include "watchdog_resen_test.sv"
	`include "watchdog_disable_inter_test.sv"
	`include "watchdog_lock_test.sv"
	`include "watchdog_PeripheralID_check_test.sv"
	
`endif  //WATCHDOG_TEST_SVH
