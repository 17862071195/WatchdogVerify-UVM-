class c_6_3;
    rand integer delay; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq_lib/watchdog_resen_virtual_sequence.sv:21)
    {
       (delay inside {[5:3]});
    }
endclass

program p_6_3;
    c_6_3 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xz1zzxzx0zzxxzzz0zz1z1xz11zzz0xxxzxxzxxxzxzzzxzxzzzxxxxxzxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
