`ifndef WATCHDOG_COVERAGE_SVH
`define WATCHDOG_COVERAGE_SVH

	`include "watchdog_coverage_module.sv"

`endif