`ifndef WATCHDOG_CONFIG_SVH
`define WATCHDOG_CONFIG_SVH

  `include "watchdog_config.sv"


`endif  //WATCHDOG_FONFIG_SVH