`ifndef WATCHDOG_REG_SVH
`define WATCHDOG_REG_SVH

	`include "watchdog_reg.sv"

`endif