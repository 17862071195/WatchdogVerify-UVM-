class c_49_3;
    rand integer delay; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq_lib/watchdog_resen_virtual_sequence.sv:21)
    {
       (delay inside {[5:3]});
    }
endclass

program p_49_3;
    c_49_3 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11x1z1111z01z100010zzzzx11z0011xzxxxxzxxxxxzzzzxxzxxxxzzxxxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
